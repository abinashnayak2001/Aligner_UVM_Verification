///////////////////////////////////////////////////////////////////////////////
// File:        cfs_algn_test_defines.sv
// Author:      Cristian Florin Slav
// Date:        2023-12-02
// Description: Defines required by the Aligner tests.
///////////////////////////////////////////////////////////////////////////////
`ifndef CFS_ALGN_TEST_DEFINES_SV
  `define CFS_ALGN_TEST_DEFINES_SV

  `ifndef CFS_ALGN_TEST_ALGN_DATA_WIDTH
    `define CFS_ALGN_TEST_ALGN_DATA_WIDTH 32
  `endif

`endif
